package init_fifo

import FIFOF::*;
import RegFile::*;

module mkInitFifo(Empty);
	
	

endmodule


endpackage